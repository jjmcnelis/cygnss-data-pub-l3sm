netcdf _ucar_cu_cygnss_sm_v1_2018_122 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 252 ;
	lon = 802 ;
	timeslices = 4 ;
	startstop = 2 ;
variables:
	float time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:units = "days since 1970-01-01 00:00:00 UTC" ;
		time:coverage_content_type = "coordinate" ;
	float latitude(lon, lat) ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "latitude" ;
		latitude:axis = "Y" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "coordinate" ;
	float longitude(lon, lat) ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "longitude" ;
		longitude:axis = "X" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "coordinate" ;
	float timeintervals(startstop, timeslices) ;
		timeintervals:long_name = "start and stop time for the sub-daily time periods" ;
		timeintervals:units = "hours" ;
		timeintervals:coverage_content_type = "referenceInformation" ;
	float SIGMA_daily(lon, lat) ;
		SIGMA_daily:_FillValue = -9999.f ;
		SIGMA_daily:comment = "units represent soil moisture content as a fractional volume (cm3 cm-3)" ;
		SIGMA_daily:long_name = "standard deviation of soil moisture retrievals during the 24 hr period for the grid cell" ;
		SIGMA_daily:units = "1" ;
		SIGMA_daily:coverage_content_type = "modelResult" ;
	float SM_daily(lon, lat) ;
		SM_daily:_FillValue = -9999.f ;
		SM_daily:comment = "units represent soil moisture content as a fractional volume (cm3 cm-3)" ;
		SM_daily:long_name = "mean soil moisture retrieval during the daily time periods for the grid cell" ;
		SM_daily:units = "1" ;
		SM_daily:coverage_content_type = "modelResult" ;
	float SM_subdaily(timeslices, lon, lat) ;
		SM_subdaily:_FillValue = -9999.f ;
		SM_subdaily:comment = "units represent soil moisture content as a fractional volume (cm3 cm-3)" ;
		SM_subdaily:long_name = "mean soil moisture retrieval during the sub-daily time periods for the grid cell" ;
		SM_subdaily:units = "1" ;
		SM_subdaily:coverage_content_type = "modelResult" ;
	float SIGMA_subdaily(timeslices, lon, lat) ;
		SIGMA_subdaily:_FillValue = -9999.f ;
		SIGMA_subdaily:comment = "units represent soil moisture content as a fractional volume (cm3 cm-3)" ;
		SIGMA_subdaily:long_name = "standard deviation of soil moisture retrievals during the sub-daily time periods for the grid cell" ;
		SIGMA_subdaily:units = "1" ;
		SIGMA_subdaily:coverage_content_type = "modelResult" ;

// global attributes:
		:source = "ucar_cu_cygnss_sm_v1_2018_122.nc" ;
		:id = "PODAAC-CYGNS-L3SM1" ;
		:ShortName = "CYGNSS_L3_SOIL_MOISTURE_V1.0" ;
		:title = "UCAR/CU CYGNSS Level 3 Soil Moisture Product" ;
		string :summary = "The UCAR/CU Cyclone Global Navigation Satellite System (CYGNSS) Level 3 Soil Moisture Product is an L-band bistatic radar dataset that provides estimates of 0-5 cm soil moisture at a 6-hour discretization for the majority of the extratropics. CYGNSS is a constellation of eight small satellites designed to observe ocean surface wind speed during hurricanes (PI Chris Ruf, University of Michigan); it is a NASA Earth Ventures Mission that was launched in December of 2016. These satellites employ a relatively new remote sensing technique called GNSS-Reflectometry (GNSS-R), which records L-band signals transmitted by navigation satellites that have reflected off of the Earth’s surface and back into space. Soil moisture estimates were produced by calculating the slope of the best-fit linear regression between SMAP soil moisture and CYGNSS \'effective reflectivity\', which gives reflectivity corrected for antenna gain, range, and GPS transmit power." ;
		:comment = "Dataset created by UCAR and CU Boulder" ;
		:program = "CYGNSS" ;
		:project = "CYGNSS" ;
		:institution = "COSMIC Data Analysis and Archive Center, Constellation Observing System for Meteorology, Ionosphere and Climate, University Corporation for Atmospheric Research (UCAR/COSMIC/CDAAC)" ;
		:references = "Chew, C.; Small, E. Description of the UCAR/CU Soil Moisture Product. Remote Sens. 2020, 12, 1558. https://doi.org/10.3390/rs12101558" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:keywords = "EARTH SCIENCE > LAND SURFACE > SOILS > SOIL MOISTURE/WATER CONTENT" ;
		:Conventions = "CF-1.6,ACDD-1.3" ;
		:license = "Freely Distributed" ;
		:version = 1. ;
		:history = "Created 24-Apr-2019 10:49:01Modified for PODAAC release 2020-09-24T04:02:54" ;
		:cdm_data_type = "Grid" ;
		:creator_name = "Clara Chew, Eric Small" ;
		:creator_type = "person, person" ;
		:creator_url = "https://staff.ucar.edu/users/clarac, http://geode.colorado.edu/~small/" ;
		:creator_email = "claraac@ucar.edu, eric.small@colorado.edu" ;
		:creator_institution = "UCAR/COSMIC/CDAAC, UCO" ;
		:publisher_name = "PO.DAAC" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:processing_level = "3" ;
		:geospatial_lat_min = -38.14157f ;
		:geospatial_lat_max = 38.14157f ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_min = -135.f ;
		:geospatial_lon_max = 164.1286f ;
		:geospatial_lon_units = "degrees_east" ;
		:time_coverage_start = "2018-05-02T00:00:00" ;
		:time_coverage_end = "2018-05-02T23:59:59" ;
		:time_coverage_duration = "P1D" ;
		:date_created = "2019-04-24T00:00:00" ;
		:date_modified = "2020-09-24T04:02:54" ;
		:date_issued = "2020-09-24T04:02:54" ;
}

netcdf _ucar_cu_cygnss_sm_v1_static_flags {
dimensions:
	lat = 252 ;
	lon = 802 ;
variables:
	float latitude(lon, lat) ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "latitude" ;
		latitude:axis = "Y" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "coordinate" ;
	float longitude(lon, lat) ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "longitude" ;
		longitude:axis = "X" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "coordinate" ;
	ubyte flag_small_SM_range(lon, lat) ;
		flag_small_SM_range:long_name = "Small data range flag" ;
		flag_small_SM_range:comment = "Indicates that CYGNSS was calibrated to SMAP data with a small range of soil moisture values (< 0.1 cm3 cm-3), which means the uncertainty in beta is large." ;
		flag_small_SM_range:valid_range = 0UB, 1UB ;
		flag_small_SM_range:flag_values = 0UB, 1UB ;
		flag_small_SM_range:flag_meanings = "normal_range small_range" ;
	ubyte flag_poor_SMAP(lon, lat) ;
		flag_poor_SMAP:long_name = "SMAP soil moisture retrieval quality flag" ;
		flag_poor_SMAP:comment = "Indicates that CYGNSS was calibrated to SMAP data where a large portion (>90%) of the SMAP soil moisture retrievals were flagged as ‘not recommended for retrieval.’" ;
		flag_poor_SMAP:valid_range = 0UB, 1UB ;
		flag_poor_SMAP:flag_values = 0UB, 1UB ;
		flag_poor_SMAP:flag_meanings = "normal_smap_soil_moisture_quality low_smap_soil_moisture_quality" ;
	ubyte flag_high_ubrmsd(lon, lat) ;
		flag_high_ubrmsd:long_name = "High unbiased RMS difference flag" ;
		flag_high_ubrmsd:comment = "Indicates a high unbiased root mean square difference between CYGNSS and SMAP retrievals (> 0.08 cm3 cm-3)." ;
		flag_high_ubrmsd:valid_range = 0UB, 1UB ;
		flag_high_ubrmsd:flag_values = 0UB, 1UB ;
		flag_high_ubrmsd:flag_meanings = "normal_unbiased_rms_difference high_unbiased_rms_difference" ;
	ubyte flag_few_obs(lon, lat) ;
		flag_few_obs:long_name = "Low observation count flag" ;
		flag_few_obs:comment = "Indicates a small number of observations in the grid cell for calibration, leading to a less certain beta (n < 100)." ;
		flag_few_obs:valid_range = 0UB, 1UB ;
		flag_few_obs:flag_values = 0UB, 1UB ;
		flag_few_obs:flag_meanings = "normal_number_of_calibration_observations low_number_of_calibration_observations" ;
	ubyte flag_low_signal(lon, lat) ;
		flag_low_signal:long_name = "Low mean effective reflectivity flag" ;
		flag_low_signal:comment = "Indicates low mean Pr,eff after water point removal in the cell, which likely means that roughness or vegetation effects are dominate (mean Pr,eff < 5 dB)." ;
		flag_low_signal:valid_range = 0UB, 1UB ;
		flag_low_signal:flag_values = 0UB, 1UB ;
		flag_low_signal:flag_meanings = "normal_mean_preff low_mean_preff" ;

// global attributes:
		:source = "ucar_cu_cygnss_sm_v1_static_flags.nc" ;
		:id = "PODAAC-CYGNU-L3SM1" ;
		:ShortName = "CYGNSS_L3_SOIL_MOISTURE_V1.0" ;
		:title = "UCAR/CU CYGNSS Level 3 Soil Moisture Product" ;
		:summary = "CYGNSS soil moisture static quality flag file" ;
		:comment = "Dataset created by UCAR and CU Boulder" ;
		:program = "CYGNSS" ;
		:project = "CYGNSS" ;
		:institution = "COSMIC Data Analysis and Archive Center, Constellation Observing System for Meteorology, Ionosphere and Climate, University Corporation for Atmospheric Research (UCAR/COSMIC/CDAAC)" ;
		:references = "Chew, C.; Small, E. Description of the UCAR/CU Soil Moisture Product. Remote Sens. 2020, 12, 1558. https://doi.org/10.3390/rs12101558" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:keywords = "EARTH SCIENCE > LAND SURFACE > SOILS > SOIL MOISTURE/WATER CONTENT" ;
		:Conventions = "CF-1.6,ACDD-1.3" ;
		:license = "Freely Distributed" ;
		:version = 1. ;
		:history = "Created 24-Apr-2019 10:48:14. Modified for PODAAC release 2020-10-13T22:25:30." ;
		:cdm_data_type = "Grid" ;
		:creator_name = "Clara Chew, Eric Small" ;
		:creator_type = "person, person" ;
		:creator_url = "https://staff.ucar.edu/users/clarac, http://geode.colorado.edu/~small/" ;
		:creator_email = "claraac@ucar.edu, eric.small@colorado.edu" ;
		:creator_institution = "UCAR/COSMIC/CDAAC, UCO" ;
		:publisher_name = "PO.DAAC" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:processing_level = "3" ;
		:geospatial_lat_min = -38.14157f ;
		:geospatial_lat_max = 38.14157f ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_min = -135.f ;
		:geospatial_lon_max = 164.1286f ;
		:geospatial_lon_units = "degrees_east" ;
		:date_created = "2019-04-24T00:00:00" ;
		:date_modified = "2020-10-13T22:25:30" ;
		:date_issued = "2020-10-13T22:25:30" ;
}

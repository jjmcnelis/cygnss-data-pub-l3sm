netcdf _ucar_cu_cygnss_sm_v1_2020_134 {
dimensions:
	time = 1 ;
	lat = 252 ;
	lon = 802 ;
	timeslices = 4 ;
	startstop = 2 ;
variables:
	float time(time) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "days since 1970-01-01 00:00:00 UTC" ;
		time:coverage_content_type = "referenceInformation" ;
	float latitude(lat, lon) ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "latitude" ;
		latitude:axis = "Y" ;
		latitude:units = "degrees_north" ;
		latitude:coverage_content_type = "coordinate" ;
	float longitude(lat, lon) ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "longitude" ;
		longitude:axis = "X" ;
		longitude:units = "degrees_east" ;
		longitude:coverage_content_type = "coordinate" ;
	float SM_daily(time, lat, lon) ;
		SM_daily:_FillValue = -9999.f ;
		SM_daily:comment = "units represent soil moisture content as a fractional volume (cm3 cm-3)" ;
		SM_daily:long_name = "mean soil moisture retrieval during the daily time periods for the grid cell" ;
		SM_daily:units = "1" ;
		SM_daily:coverage_content_type = "modelResult" ;
	float SM_subdaily(timeslices, lat, lon) ;
		SM_subdaily:_FillValue = -9999.f ;
		SM_subdaily:comment = "units represent soil moisture content as a fractional volume (cm3 cm-3)" ;
		SM_subdaily:long_name = "mean soil moisture retrieval during the sub-daily time periods for the grid cell" ;
		SM_subdaily:units = "1" ;
		SM_subdaily:coverage_content_type = "modelResult" ;
	float SIGMA_daily(time, lat, lon) ;
		SIGMA_daily:_FillValue = -9999.f ;
		SIGMA_daily:comment = "units represent soil moisture content as a fractional volume (cm3 cm-3)" ;
		SIGMA_daily:long_name = "standard deviation of soil moisture retrievals during the 24 hr period for the grid cell" ;
		SIGMA_daily:units = "1" ;
		SIGMA_daily:coverage_content_type = "modelResult" ;
	float SIGMA_subdaily(timeslices, lat, lon) ;
		SIGMA_subdaily:_FillValue = -9999.f ;
		SIGMA_subdaily:comment = "units represent soil moisture content as a fractional volume (cm3 cm-3)" ;
		SIGMA_subdaily:long_name = "standard deviation of soil moisture retrievals during the sub-daily time periods for the grid cell" ;
		SIGMA_subdaily:units = "1" ;
		SIGMA_subdaily:coverage_content_type = "modelResult" ;
	float timeintervals(timeslices, startstop) ;
		timeintervals:_FillValue = -9999.f ;
		timeintervals:long_name = "start and stop time for the sub-daily time periods" ;
		timeintervals:units = "hours" ;
		timeintervals:coverage_content_type = "referenceInformation" ;

// global attributes:
		:source = "ucar_cu_cygnss_sm_v1_2020_134.nc" ;
		:id = "PODAAC-CYGNU-L3SM1" ;
		:ShortName = "CYGNSS_L3_SOIL_MOISTURE_V1.0" ;
		:title = "CYGNSS Level 3 Soil Moisture from UCAR/CU" ;
		:summary = "The CYGNSS Level 3 Soil Moisture Product provides volumetric water content estimates for soils between 0-5 cm depth at a 6-hour discretization for most of the subtropics. The data were produced by CYGNSS investigators at the University Corporation for Atmospheric Research (UCAR) and the University Colorado at Boulder (CU), and derive from version 2.1 of the CYGNSS L1 SDR. The soil moisture algorithm uses collocated soil moisture retrievals from SMAP to calibrate CYGNSS observations from the same day. For a given location, a linear relationship between the SMAP soil moisture and CYGNSS reflectivity is determined and used to transform the CYGNSS observations into soil moisture. The data are archived in daily files in netCDF-4 format. Two soil moisture variables report the volumetric water content in units of cm3/cm3. The variable SM_subdaily includes up to four soil moisture estimates per day. Another variable SM_daily provides a daily average. The time series covers the period from March 2017 to August 2020." ;
		:comment = "Dataset created by UCAR and CU Boulder" ;
		:program = "CYGNSS" ;
		:project = "CYGNSS" ;
		:institution = "COSMIC Data Analysis and Archive Center, Constellation Observing System for Meteorology, Ionosphere and Climate, University Corporation for Atmospheric Research (UCAR/COSMIC/CDAAC)" ;
		:references = "Chew, C.; Small, E. Description of the UCAR/CU Soil Moisture Product. Remote Sens. 2020, 12, 1558. https://doi.org/10.3390/rs12101558" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:keywords = "EARTH SCIENCE > LAND SURFACE > SOILS > SOIL MOISTURE/WATER CONTENT" ;
		:Conventions = "CF-1.6,ACDD-1.3" ;
		:license = "Freely Distributed" ;
		:version = 1. ;
		:history = "Created 2020-05-28 02:28:59.624705. Modified for PODAAC release 2020-10-31T02:08:56." ;
		:cdm_data_type = "Grid" ;
		:creator_name = "Clara Chew, Eric Small" ;
		:creator_type = "person, person" ;
		:creator_url = "https://staff.ucar.edu/users/clarac, http://geode.colorado.edu/~small/" ;
		:creator_email = "claraac@ucar.edu, eric.small@colorado.edu" ;
		:creator_institution = "UCAR/COSMIC/CDAAC, UCO" ;
		:publisher_name = "PO.DAAC" ;
		:publisher_email = "podaac@podaac.jpl.nasa.gov" ;
		:publisher_type = "institution" ;
		:publisher_url = "https://podaac.jpl.nasa.gov" ;
		:publisher_institution = "NASA/JPL/PODAAC" ;
		:processing_level = "3" ;
		:geospatial_lat_min = -38.14157f ;
		:geospatial_lat_max = 38.14157f ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_min = -135.f ;
		:geospatial_lon_max = 164.1286f ;
		:geospatial_lon_units = "degrees_east" ;
		:time_coverage_start = "2020-05-13T00:00:00" ;
		:time_coverage_end = "2020-05-13T23:59:59" ;
		:time_coverage_duration = "P1D" ;
		:date_created = "2020-05-28T00:00:00" ;
		:date_modified = "2020-10-31T02:08:56" ;
		:date_issued = "2020-10-31T02:08:56" ;
}
